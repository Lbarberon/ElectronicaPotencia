** Profile: "SCHEMATIC1-CargaRL"  [ C:\Users\lucho\OneDrive\Escritorio\ElectronicaPotencia-main\TP3\Simulacion\tp3_ep-pspicefiles\schematic1\cargarl.sim ] 

** Creating circuit file "CargaRL.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\lucho\cdssetup\OrCAD_PSpice\23.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 80ms 40ms 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
