** Profile: "SCHEMATIC1-Carga_R"  [ C:\Users\lucho\OneDrive\Escritorio\ElectronicaPotencia-main\ElectronicaPotencia-main\ElectronicaPotencia-main\TP3\Simulacion\tp3_ep-pspicefiles\schematic1\carga_r.sim ] 

** Creating circuit file "Carga_R.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\lucho\cdssetup\OrCAD_PSpice\23.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 80m 40m 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
