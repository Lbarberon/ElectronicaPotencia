** Profile: "SCHEMATIC1-CargaRL1"  [ C:\Users\lucho\OneDrive\Escritorio\ElectronicaPotencia-main\TP3\Simulacion\TP3_EP-PSpiceFiles\SCHEMATIC1\CargaRL1.sim ] 

** Creating circuit file "CargaRL1.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\lucho\cdssetup\OrCAD_PSpice\23.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 100ms 40ms 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
